
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_top_kernel.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_top_kernel.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_top_kernel.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;

    seq_loop_intf#(4) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ST_fsm_state1;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ST_fsm_state1;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.ap_ST_fsm_state4;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(4) seq_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_54_1_fu_1154.grp_top_kernel_Pipeline_VITIS_LOOP_56_2_fu_1090.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1;
    assign upc_loop_intf_2.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_2.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_2.iter_start_enable = 1'b1;
    assign upc_loop_intf_2.iter_end_enable = 1'b1;
    assign upc_loop_intf_2.quit_enable = 1'b1;
    assign upc_loop_intf_2.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_83_6_fu_1686.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_3.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_3.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_5_fu_1747.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_4.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_4.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_51_fu_2011.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_5.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_5.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_52_fu_2275.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_6.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_6.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_53_fu_2539.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_7.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_7.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_54_fu_2803.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_8.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_8.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_55_fu_3067.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_9.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_9.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_56_fu_3331.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_10.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_enable_reg_pp0_iter44;
    assign upc_loop_intf_10.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_69_4_VITIS_LOOP_71_57_fu_3595.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_9_fu_3859.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_12.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_12.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_98_fu_3873.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_13.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_13.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_99_fu_3936.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_14.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_14.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_910_fu_3971.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_15.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_15.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_911_fu_4034.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_16.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_16.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_912_fu_4055.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_17.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_17.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_913_fu_4118.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b1;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(1) upc_loop_monitor_17;
    upc_loop_intf#(1) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_18.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_18.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_90_8_VITIS_LOOP_91_914_fu_4153.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b1;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(1) upc_loop_monitor_18;
    upc_loop_intf#(1) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_99_10_fu_4216.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b1;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(1) upc_loop_monitor_19;
    upc_loop_intf#(1) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_13_fu_4348.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b1;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(1) upc_loop_monitor_20;
    upc_loop_intf#(1) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_21.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_21.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1315_fu_4378.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b1;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(1) upc_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_22.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_22.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1316_fu_4457.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b1;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(1) upc_loop_monitor_22;
    upc_loop_intf#(1) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_23.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_23.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1317_fu_4508.ap_done_int;
    assign upc_loop_intf_23.loop_continue = 1'b1;
    assign upc_loop_intf_23.quit_at_end = 1'b1;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(1) upc_loop_monitor_23;
    upc_loop_intf#(1) upc_loop_intf_24(clock,reset);
    assign upc_loop_intf_24.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_CS_fsm;
    assign upc_loop_intf_24.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_24.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_24.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_start;
    assign upc_loop_intf_24.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_ready;
    assign upc_loop_intf_24.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1318_fu_4587.ap_done_int;
    assign upc_loop_intf_24.loop_continue = 1'b1;
    assign upc_loop_intf_24.quit_at_end = 1'b1;
    assign upc_loop_intf_24.finish = finish;
    csv_file_dump upc_loop_csv_dumper_24;
    upc_loop_monitor #(1) upc_loop_monitor_24;
    upc_loop_intf#(1) upc_loop_intf_25(clock,reset);
    assign upc_loop_intf_25.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_CS_fsm;
    assign upc_loop_intf_25.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_25.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_25.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_start;
    assign upc_loop_intf_25.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_ready;
    assign upc_loop_intf_25.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1319_fu_4624.ap_done_int;
    assign upc_loop_intf_25.loop_continue = 1'b1;
    assign upc_loop_intf_25.quit_at_end = 1'b1;
    assign upc_loop_intf_25.finish = finish;
    csv_file_dump upc_loop_csv_dumper_25;
    upc_loop_monitor #(1) upc_loop_monitor_25;
    upc_loop_intf#(1) upc_loop_intf_26(clock,reset);
    assign upc_loop_intf_26.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_CS_fsm;
    assign upc_loop_intf_26.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_26.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_26.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_26.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_start;
    assign upc_loop_intf_26.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_ready;
    assign upc_loop_intf_26.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1320_fu_4703.ap_done_int;
    assign upc_loop_intf_26.loop_continue = 1'b1;
    assign upc_loop_intf_26.quit_at_end = 1'b1;
    assign upc_loop_intf_26.finish = finish;
    csv_file_dump upc_loop_csv_dumper_26;
    upc_loop_monitor #(1) upc_loop_monitor_26;
    upc_loop_intf#(1) upc_loop_intf_27(clock,reset);
    assign upc_loop_intf_27.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_CS_fsm;
    assign upc_loop_intf_27.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_27.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_27.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_start;
    assign upc_loop_intf_27.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_ready;
    assign upc_loop_intf_27.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_12_VITIS_LOOP_110_1321_fu_4754.ap_done_int;
    assign upc_loop_intf_27.loop_continue = 1'b1;
    assign upc_loop_intf_27.quit_at_end = 1'b1;
    assign upc_loop_intf_27.finish = finish;
    csv_file_dump upc_loop_csv_dumper_27;
    upc_loop_monitor #(1) upc_loop_monitor_27;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);
    upc_loop_csv_dumper_24 = new("./upc_loop_status24.csv");
    upc_loop_monitor_24 = new(upc_loop_intf_24,upc_loop_csv_dumper_24);
    upc_loop_csv_dumper_25 = new("./upc_loop_status25.csv");
    upc_loop_monitor_25 = new(upc_loop_intf_25,upc_loop_csv_dumper_25);
    upc_loop_csv_dumper_26 = new("./upc_loop_status26.csv");
    upc_loop_monitor_26 = new(upc_loop_intf_26,upc_loop_csv_dumper_26);
    upc_loop_csv_dumper_27 = new("./upc_loop_status27.csv");
    upc_loop_monitor_27 = new(upc_loop_intf_27,upc_loop_csv_dumper_27);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_24);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_26);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_27);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
